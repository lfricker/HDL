//---------------------------------
// Projet : HDL_2020
// Name   : memory
// Author : lfr
// Date   : 14.01.2021
//---------------------------------


module memory
(

);



endmodule